module Hello;
 initial begin $display("Hello World"); $finish; end
endmodule